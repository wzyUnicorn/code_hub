class vseq_lpc_beep extends uvm_sequence;
    `uvm_object_utils(vseq_lpc_beep)
    `uvm_declare_p_sequencer(virtual_sequencer)

    virtual task body();
        btn_base_sequence btn_seq;
        lpc_transaction tr;

    if(starting_phase!=null) starting_phase.raise_objection(this);
        `uvm_do_on(btn_seq,p_sequencer.vbtn_sqr) // button power on
    for(int i=0;i<5;i++) begin
        // lpc control buzzer frequency
        `uvm_do_on_with(tr,p_sequencer.vlpc_sqr,{tr.cyctype==4'b0010;tr.addr==16'h0808;tr.dataIn=={5'b00001<<i,3'b001};})
    end
    if(starting_phase!=null) starting_phase.drop_objection(this);
    endtask
endclass
