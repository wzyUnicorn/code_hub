interface cnn_if;
    logic cnn_done_irq;
endinterface: cnn_if
