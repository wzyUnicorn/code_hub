package test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import btn_agent_pkg::*;
    import iic_agent_pkg::*;
    import lpc_agent_pkg::*;
    import tele_agent_pkg::*;
    import env_pkg::*;

    `include "virtual_sequencer.sv"
    `include "seqlib/virtual_sequence_base.sv"
    `include "seqlib/vseq_btn_power_on_off.sv"
    `include "seqlib/vseq_btn_power_on_reset.sv"
    `include "seqlib/vseq_btn_power_on_interrupt.sv"
    `include "seqlib/vseq_btn_power_on_dcok.sv"
    `include "seqlib/vseq_btn_power_on_alarm.sv"
    `include "seqlib/vseq_btn_power_on_jitter.sv"
    `include "seqlib/vseq_btn_power_on_again.sv"
    `include "seqlib/vseq_iic_power_on_off.sv"
    `include "seqlib/vseq_iic_power_on_reset.sv"
    `include "seqlib/vseq_iic_power_on_mtrst.sv"
    `include "seqlib/vseq_iic_power_on_beep.sv"
    `include "seqlib/vseq_lpc_power_off.sv"
    `include "seqlib/vseq_lpc_vga.sv"
    `include "seqlib/vseq_lpc_vga_disable.sv"
    `include "seqlib/vseq_lpc_soft_reset.sv"
    `include "seqlib/vseq_lpc_mt_reset.sv"
    `include "seqlib/vseq_lpc_ich.sv"
    `include "seqlib/vseq_lpc_beep.sv"
    `include "seqlib/vseq_lpc_write_read.sv"
    `include "seqlib/vseq_lpc_transfer_abort.sv"
    `include "seqlib/vseq_btn_on_iic_reset.sv"
    `include "seqlib/vseq_btn_on_iic_off.sv"
    `include "seqlib/vseq_btn_on_iic_beep.sv"
    `include "seqlib/vseq_btn_on_iic_random_addr.sv"
    `include "seqlib/vseq_btn_on_tele_off.sv"
    `include "seqlib/vseq_btn_on_tele_reset.sv"
    `include "seqlib/vseq_iic_on_btn_reset.sv"
    `include "seqlib/vseq_iic_on_btn_off.sv"
    `include "seqlib/vseq_iic_on_lpc_reset.sv"
    `include "seqlib/vseq_iic_on_lpc_mtrst.sv"
    `include "seqlib/vseq_iic_on_lpc_off.sv"
    `include "seqlib/vseq_iic_on_lpc_vga.sv"
    `include "seqlib/vseq_iic_on_lpc_ich.sv"
    `include "seqlib/vseq_iic_on_lpc_beep.sv"
    `include "seqlib/vseq_iic_on_tele_reset.sv"
    `include "seqlib/vseq_iic_on_tele_off.sv"
    `include "seqlib/vseq_tele_on_off.sv"
    `include "seqlib/vseq_tele_on_rst_off.sv"
    `include "seqlib/vseq_tele_on_btn_off.sv"
    `include "seqlib/vseq_tele_on_btn_reset.sv"
    `include "seqlib/vseq_tele_on_iic_reset.sv"
    `include "seqlib/vseq_tele_on_iic_off.sv"
    `include "seqlib/vseq_tele_on_lpc_reset.sv"
    `include "seqlib/vseq_tele_on_lpc_off.sv"

    `include "test_base.sv"
    `include "test_btn_power_on_off.sv"
    `include "test_btn_power_on_reset.sv"
    `include "test_btn_power_on_interrupt.sv"
    `include "test_btn_power_on_dcok.sv"
    `include "test_btn_power_on_alarm.sv"
    `include "test_btn_power_on_jitter.sv"
    `include "test_btn_power_on_again.sv"
    `include "test_iic_power_on_off.sv"
    `include "test_iic_power_on_reset.sv"
    `include "test_iic_power_on_mtrst.sv"
    `include "test_iic_power_on_beep.sv"
    `include "test_lpc_power_off.sv"
    `include "test_lpc_soft_reset.sv"
    `include "test_lpc_mt_reset.sv"
    `include "test_lpc_vga.sv"
    `include "test_lpc_vga_disable.sv"
    `include "test_lpc_ich.sv"
    `include "test_lpc_beep.sv"
    `include "test_lpc_write_read.sv"
    `include "test_lpc_transfer_abort.sv"
    `include "test_btn_on_iic_reset.sv"
    `include "test_btn_on_iic_off.sv"
    `include "test_btn_on_iic_beep.sv"
    `include "test_btn_on_iic_random_addr.sv"
    `include "test_btn_on_tele_off.sv"
    `include "test_btn_on_tele_reset.sv"
    `include "test_iic_on_btn_reset.sv"
    `include "test_iic_on_btn_off.sv"
    `include "test_iic_on_lpc_reset.sv"
    `include "test_iic_on_lpc_mtrst.sv"
    `include "test_iic_on_lpc_off.sv"
    `include "test_iic_on_lpc_vga.sv"
    `include "test_iic_on_lpc_ich.sv"
    `include "test_iic_on_lpc_beep.sv"
    `include "test_iic_on_tele_reset.sv"
    `include "test_iic_on_tele_off.sv"
    `include "test_tele_on_off.sv"
    `include "test_tele_on_rst_off.sv"
    `include "test_tele_on_btn_off.sv"
    `include "test_tele_on_btn_reset.sv"
    `include "test_tele_on_iic_reset.sv"
    `include "test_tele_on_iic_off.sv"
    `include "test_tele_on_lpc_reset.sv"
    `include "test_tele_on_lpc_off.sv"
endpackage
