/**********************************
copyright@FPGA OPEN SOURCE STUDIO
微信公众号：FPGA开源工作室
***********************************/
`timescale 1ns / 1ps

module rom_sw(
input  clk,
input [8:0] addr,
output signed [31:0] dout);
(*rom_style = "block" *) reg signed [31:0] data;
always @(posedge clk) 
begin
    case(addr)
      0:data<=32'd0;
      1:data<=32'd485243364;
      2:data<=32'd894802018;
      3:data<=32'd1191737781;
      4:data<=32'd1352751513;
      5:data<=32'd1370062590;
      6:data<=32'd1251556367;
      7:data<=32'd1019232785;
      8:data<=32'd706170578;
      9:data<=32'd352376348;
      10:data<=32'd0;
      11:data<=-32'd311543726;
      12:data<=-32'd550009086;
      13:data<=-32'd693829686;
      14:data<=-32'd734336548;
      15:data<=-32'd676457349;
      16:data<=-32'd537793542;
      17:data<=-32'd345767722;
      18:data<=-32'd126503314;
      19:data<=32'd0;
      20:data<=32'd0;
      21:data<=32'd0;
      22:data<=32'd0;
      23:data<=32'd0;
      24:data<=32'd0;
      25:data<=32'd0;
      26:data<=32'd0;
      27:data<=32'd0;
      28:data<=32'd0;
      29:data<=32'd0;
      30:data<=32'd0;
      31:data<=32'd0;
      32:data<=32'd0;
      33:data<=32'd0;
      34:data<=32'd0;
      35:data<=32'd0;
      36:data<=32'd0;
      37:data<=32'd0;
      38:data<=32'd0;
      39:data<=32'd0;
      40:data<=32'd0;
      41:data<=32'd0;
      42:data<=32'd0;
      43:data<=32'd0;
      44:data<=32'd0;
      45:data<=32'd0;
      46:data<=32'd0;
      47:data<=32'd0;
      48:data<=32'd0;
      49:data<=32'd0;
      50:data<=32'd0;
      51:data<=32'd0;
      52:data<=32'd0;
      53:data<=32'd0;
      54:data<=32'd0;
      55:data<=32'd0;
      56:data<=32'd0;
      57:data<=32'd0;
      58:data<=32'd0;
      59:data<=32'd0;
      60:data<=32'd0;
      61:data<=32'd0;
      62:data<=32'd0;
      63:data<=32'd0;
      64:data<=32'd0;
      65:data<=32'd0;
      66:data<=32'd0;
      67:data<=32'd0;
      68:data<=32'd0;
      69:data<=32'd0;
      70:data<=32'd0;
      71:data<=32'd0;
      72:data<=32'd0;
      73:data<=32'd0;
      74:data<=32'd0;
      75:data<=32'd0;
      76:data<=32'd0;
      77:data<=32'd0;
      78:data<=32'd0;
      79:data<=32'd0;
      80:data<=32'd0;
      81:data<=32'd0;
      82:data<=32'd0;
      83:data<=32'd0;
      84:data<=32'd0;
      85:data<=32'd0;
      86:data<=32'd0;
      87:data<=32'd0;
      88:data<=32'd0;
      89:data<=32'd0;
      90:data<=32'd0;
      91:data<=32'd0;
      92:data<=32'd0;
      93:data<=32'd0;
      94:data<=32'd0;
      95:data<=32'd0;
      96:data<=32'd0;
      97:data<=32'd0;
      98:data<=32'd0;
      99:data<=32'd0;
      100:data<=32'd0;
      101:data<=32'd0;
      102:data<=32'd0;
      103:data<=32'd0;
      104:data<=32'd0;
      105:data<=32'd0;
      106:data<=32'd0;
      107:data<=32'd0;
      108:data<=32'd0;
      109:data<=32'd0;
      110:data<=32'd0;
      111:data<=32'd0;
      112:data<=32'd0;
      113:data<=32'd0;
      114:data<=32'd0;
      115:data<=32'd0;
      116:data<=32'd0;
      117:data<=32'd0;
      118:data<=32'd0;
      119:data<=32'd0;
      120:data<=32'd0;
      121:data<=32'd0;
      122:data<=32'd0;
      123:data<=32'd0;
      124:data<=32'd0;
      125:data<=32'd0;
      126:data<=32'd0;
      127:data<=32'd0;
      128:data<=32'd0;
      129:data<=32'd0;
      130:data<=32'd0;
      131:data<=32'd0;
      132:data<=32'd0;
      133:data<=32'd0;
      134:data<=32'd0;
      135:data<=32'd0;
      136:data<=32'd0;
      137:data<=32'd0;
      138:data<=32'd0;
      139:data<=32'd0;
      140:data<=32'd0;
      141:data<=32'd0;
      142:data<=32'd0;
      143:data<=32'd0;
      144:data<=32'd0;
      145:data<=32'd0;
      146:data<=32'd0;
      147:data<=32'd0;
      148:data<=32'd0;
      149:data<=32'd0;
      150:data<=32'd0;
      151:data<=32'd0;
      152:data<=32'd0;
      153:data<=32'd0;
      154:data<=32'd0;
      155:data<=32'd0;
      156:data<=32'd0;
      157:data<=32'd0;
      158:data<=32'd0;
      159:data<=32'd0;
      160:data<=32'd0;
      161:data<=32'd0;
      162:data<=32'd0;
      163:data<=32'd0;
      164:data<=32'd0;
      165:data<=32'd0;
      166:data<=32'd0;
      167:data<=32'd0;
      168:data<=32'd0;
      169:data<=32'd0;
      170:data<=32'd0;
      171:data<=32'd0;
      172:data<=32'd0;
      173:data<=32'd0;
      174:data<=32'd0;
      175:data<=32'd0;
      176:data<=32'd0;
      177:data<=32'd0;
      178:data<=32'd0;
      179:data<=32'd0;
      180:data<=32'd0;
      181:data<=32'd0;
      182:data<=32'd0;
      183:data<=32'd0;
      184:data<=32'd0;
      185:data<=32'd0;
      186:data<=32'd0;
      187:data<=32'd0;
      188:data<=32'd0;
      189:data<=32'd0;
      190:data<=32'd0;
      191:data<=32'd0;
      192:data<=32'd0;
      193:data<=32'd0;
      194:data<=32'd0;
      195:data<=32'd0;
      196:data<=32'd0;
      197:data<=32'd0;
      198:data<=32'd0;
      199:data<=32'd0;
      200:data<=32'd0;
      201:data<=32'd0;
      202:data<=32'd0;
      203:data<=32'd0;
      204:data<=32'd0;
      205:data<=32'd0;
      206:data<=32'd0;
      207:data<=32'd0;
      208:data<=32'd0;
      209:data<=32'd0;
      210:data<=32'd0;
      211:data<=32'd0;
      212:data<=32'd0;
      213:data<=32'd0;
      214:data<=32'd0;
      215:data<=32'd0;
      216:data<=32'd0;
      217:data<=32'd0;
      218:data<=32'd0;
      219:data<=32'd0;
      220:data<=32'd0;
      221:data<=32'd0;
      222:data<=32'd0;
      223:data<=32'd0;
      224:data<=32'd0;
      225:data<=32'd0;
      226:data<=32'd0;
      227:data<=32'd0;
      228:data<=32'd0;
      229:data<=32'd0;
      230:data<=32'd0;
      231:data<=32'd0;
      232:data<=32'd0;
      233:data<=32'd0;
      234:data<=32'd0;
      235:data<=32'd0;
      236:data<=32'd0;
      237:data<=32'd0;
      238:data<=32'd0;
      239:data<=32'd0;
      240:data<=32'd0;
      241:data<=32'd0;
      242:data<=32'd0;
      243:data<=32'd0;
      244:data<=32'd0;
      245:data<=32'd0;
      246:data<=32'd0;
      247:data<=32'd0;
      248:data<=32'd0;
      249:data<=32'd0;
      250:data<=32'd0;
      251:data<=32'd0;
      252:data<=32'd0;
      253:data<=32'd0;
      254:data<=32'd0;
      255:data<=32'd0;
      256:data<=32'd0;
      257:data<=32'd0;
      258:data<=32'd0;
      259:data<=32'd0;
      260:data<=32'd0;
      261:data<=32'd0;
      262:data<=32'd0;
      263:data<=32'd0;
      264:data<=32'd0;
      265:data<=32'd0;
      266:data<=32'd0;
      267:data<=32'd0;
      268:data<=32'd0;
      269:data<=32'd0;
      270:data<=32'd0;
      271:data<=32'd0;
      272:data<=32'd0;
      273:data<=32'd0;
      274:data<=32'd0;
      275:data<=32'd0;
      276:data<=32'd0;
      277:data<=32'd0;
      278:data<=32'd0;
      279:data<=32'd0;
      280:data<=32'd0;
      281:data<=32'd0;
      282:data<=32'd0;
      283:data<=32'd0;
      284:data<=32'd0;
      285:data<=32'd0;
      286:data<=32'd0;
      287:data<=32'd0;
      288:data<=32'd0;
      289:data<=32'd0;
      290:data<=32'd0;
      291:data<=32'd0;
      292:data<=32'd0;
      293:data<=32'd0;
      294:data<=32'd0;
      295:data<=32'd0;
      296:data<=32'd0;
      297:data<=32'd0;
      298:data<=32'd0;
      299:data<=32'd0;
      300:data<=32'd0;
      301:data<=32'd0;
      302:data<=32'd0;
      303:data<=32'd0;
      304:data<=32'd0;
      305:data<=32'd0;
      306:data<=32'd0;
      307:data<=32'd0;
      308:data<=32'd0;
      309:data<=32'd0;
      310:data<=32'd0;
      311:data<=32'd0;
      312:data<=32'd0;
      313:data<=32'd0;
      314:data<=32'd0;
      315:data<=32'd0;
      316:data<=32'd0;
      317:data<=32'd0;
      318:data<=32'd0;
      319:data<=32'd0;
      320:data<=32'd0;
      321:data<=32'd0;
      322:data<=32'd0;
      323:data<=32'd0;
      324:data<=32'd0;
      325:data<=32'd0;
      326:data<=32'd0;
      327:data<=32'd0;
      328:data<=32'd0;
      329:data<=32'd0;
      330:data<=32'd0;
      331:data<=32'd0;
      332:data<=32'd0;
      333:data<=32'd0;
      334:data<=32'd0;
      335:data<=32'd0;
      336:data<=32'd0;
      337:data<=32'd0;
      338:data<=32'd0;
      339:data<=32'd0;
      340:data<=32'd0;
      341:data<=32'd0;
      342:data<=32'd0;
      343:data<=32'd0;
      344:data<=32'd0;
      345:data<=32'd0;
      346:data<=32'd0;
      347:data<=32'd0;
      348:data<=32'd0;
      349:data<=32'd0;
      350:data<=32'd0;
      351:data<=32'd0;
      352:data<=32'd0;
      353:data<=32'd0;
      354:data<=32'd0;
      355:data<=32'd0;
      356:data<=32'd0;
      357:data<=32'd0;
      358:data<=32'd0;
      359:data<=32'd0;
      360:data<=32'd0;
      361:data<=32'd0;
      362:data<=32'd0;
      363:data<=32'd0;
      364:data<=32'd0;
      365:data<=32'd0;
      366:data<=32'd0;
      367:data<=32'd0;
      368:data<=32'd0;
      369:data<=32'd0;
      370:data<=32'd0;
      371:data<=32'd0;
      372:data<=32'd0;
      373:data<=32'd0;
      374:data<=32'd0;
      375:data<=32'd0;
      376:data<=32'd0;
      377:data<=32'd0;
      378:data<=32'd0;
      379:data<=32'd0;
      380:data<=32'd0;
      381:data<=32'd0;
      382:data<=32'd126503314;
      383:data<=32'd345767722;
      384:data<=32'd537793542;
      385:data<=32'd676457349;
      386:data<=32'd734336548;
      387:data<=32'd693829686;
      388:data<=32'd550009086;
      389:data<=32'd311543726;
      390:data<=32'd0;
      391:data<=-32'd352376348;
      392:data<=-32'd706170578;
      393:data<=-32'd1019232785;
      394:data<=-32'd1251556367;
      395:data<=-32'd1370062590;
      396:data<=-32'd1352751513;
      397:data<=-32'd1191737781;
      398:data<=-32'd894802018;
      399:data<=-32'd485243364;
      400:data<=32'd0;
    endcase
end
assign dout =data;
endmodule
