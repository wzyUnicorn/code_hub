package lpc_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "lpc_transaction.sv"
    `include "lpc_sequencer.sv"
    `include "lpc_driver.sv"
    `include "lpc_monitor.sv"
    `include "lpc_agent.sv"
endpackage
