typedef uvm_sequencer#(ahb_txn) ahb_slave_sequencer;
