package tele_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "tele_ctrl_item.sv"
    `include "tele_sequencer.sv"
    `include "tele_driver.sv"
    `include "tele_agent.sv"
endpackage
