package btn_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "cpld_output_tr.sv"
    `include "btn_sequencer.sv"
    `include "btn_driver.sv"
    `include "btn_monitor.sv"
    `include "btn_agent.sv"
endpackage
