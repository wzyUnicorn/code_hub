typedef uvm_sequencer#(isp_txn) isp_sequencer;
