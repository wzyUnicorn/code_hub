typedef uvm_sequencer#(cnn_txn) cnn_sequencer;
