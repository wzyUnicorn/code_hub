module rom_heart(
input  clk,
input [8:0] addr,
output signed [31:0] dout);
(*rom_style = "block" *) reg signed [31:0] data;
always @(posedge clk) 
begin
    case(addr)
      0:data<=32'd1168411192;
      1:data<=32'd1162720908;
      2:data<=32'd1157021085;
      3:data<=32'd1151311657;
      4:data<=32'd1145592561;
      5:data<=32'd1139863731;
      6:data<=32'd1134125099;
      7:data<=32'd1128376598;
      8:data<=32'd1122618160;
      9:data<=32'd1116849716;
      10:data<=32'd1111071197;
      11:data<=32'd1105282530;
      12:data<=32'd1099483646;
      13:data<=32'd1093674470;
      14:data<=32'd1087854930;
      15:data<=32'd1082024952;
      16:data<=32'd1076184459;
      17:data<=32'd1070333376;
      18:data<=32'd1064471626;
      19:data<=32'd1012400427;
      20:data<=32'd1052715809;
      21:data<=32'd1139363850;
      22:data<=32'd1247119426;
      23:data<=32'd1354811781;
      24:data<=32'd1442843654;
      25:data<=32'd1494415357;
      26:data<=32'd1497202900;
      27:data<=32'd1444779407;
      28:data<=32'd1337469925;
      29:data<=32'd1182482718;
      30:data<=32'd993269035;
      31:data<=32'd788160119;
      32:data<=32'd588416132;
      33:data<=32'd415891225;
      34:data<=32'd290565759;
      35:data<=32'd228216207;
      36:data<=32'd238483229;
      37:data<=32'd323559829;
      38:data<=32'd477658238;
      39:data<=32'd687332708;
      40:data<=32'd932644335;
      41:data<=32'd1189062976;
      42:data<=32'd1429919925;
      43:data<=32'd1629162243;
      44:data<=32'd1764122219;
      45:data<=32'd1818007924;
      46:data<=32'd1781844256;
      47:data<=32'd1655646375;
      48:data<=32'd1448683857;
      49:data<=32'd1178786524;
      50:data<=32'd870742391;
      51:data<=32'd553934061;
      52:data<=32'd259442241;
      53:data<=32'd16904942;
      54:data<=-32'd148548077;
      55:data<=-32'd218967780;
      56:data<=-32'd185581982;
      57:data<=-32'd49896358;
      58:data<=32'd176230299;
      59:data<=32'd471564211;
      60:data<=32'd807448232;
      61:data<=32'd1150545976;
      62:data<=32'd1466113402;
      63:data<=32'd1721474492;
      64:data<=32'd1889351551;
      65:data<=32'd1950709754;
      66:data<=32'd1896819567;
      67:data<=32'd1730315417;
      68:data<=32'd1465127397;
      69:data<=32'd1125275070;
      70:data<=32'd742627451;
      71:data<=32'd353839231;
      72:data<=-32'd3240476;
      73:data<=-32'd293333248;
      74:data<=-32'd487294285;
      75:data<=-32'd565112434;
      76:data<=-32'd518038437;
      77:data<=-32'd349616185;
      78:data<=-32'd75499098;
      79:data<=32'd277945704;
      80:data<=32'd676121139;
      81:data<=32'd1079536887;
      82:data<=32'd1447675905;
      83:data<=32'd1743010710;
      84:data<=32'd1934770055;
      85:data<=32'd2002077087;
      86:data<=32'd1936138745;
      87:data<=32'd1741257466;
      88:data<=32'd1434551487;
      89:data<=32'd1044397738;
      90:data<=32'd607738959;
      91:data<=32'd166511400;
      92:data<=-32'd236460327;
      93:data<=-32'd561698149;
      94:data<=-32'd777015327;
      95:data<=-32'd860776184;
      96:data<=-32'd804140359;
      97:data<=-32'd612059195;
      98:data<=-32'd302913941;
      99:data<=32'd93180464;
      100:data<=32'd537249431;
      101:data<=32'd985235556;
      102:data<=32'd1392311279;
      103:data<=32'd1717304137;
      104:data<=32'd1926796795;
      105:data<=32'd1998492840;
      106:data<=32'd1923509003;
      107:data<=32'd1707358368;
      108:data<=32'd1369517190;
      109:data<=32'd941607597;
      110:data<=32'd464365906;
      111:data<=-32'd16312173;
      112:data<=-32'd453864599;
      113:data<=-32'd805653550;
      114:data<=-32'd1037200004;
      115:data<=-32'd1125641116;
      116:data<=-32'd1062063353;
      117:data<=-32'd852473384;
      118:data<=-32'd517302037;
      119:data<=-32'd89481123;
      120:data<=32'd388725618;
      121:data<=32'd869831910;
      122:data<=32'd1305778289;
      123:data<=32'd1652665347;
      124:data<=32'd1875103887;
      125:data<=32'd1949750285;
      126:data<=32'd1867673479;
      127:data<=32'd1635313579;
      128:data<=32'd1273929938;
      129:data<=32'd817585243;
      130:data<=32'd309857015;
      131:data<=-32'd200405462;
      132:data<=-32'd663864903;
      133:data<=-32'd1035551243;
      134:data<=-32'd1279309772;
      135:data<=-32'd1371401596;
      136:data<=-32'd1302897512;
      137:data<=-32'd1080623795;
      138:data<=-32'd726560266;
      139:data<=-32'd275743268;
      140:data<=32'd227126130;
      141:data<=32'd732039788;
      142:data<=32'd1188580528;
      143:data<=32'd1550880068;
      144:data<=32'd1782148578;
      145:data<=32'd1858327962;
      146:data<=32'd1770505687;
      147:data<=32'd1525846810;
      148:data<=32'd1146947062;
      149:data<=32'd669665144;
      150:data<=32'd139642436;
      151:data<=-32'd392151598;
      152:data<=-32'd874412918;
      153:data<=-32'd1260545428;
      154:data<=-32'd1513256254;
      155:data<=-32'd1608250030;
      156:data<=-32'd1536655848;
      157:data<=-32'd1305944279;
      158:data<=-32'd939239885;
      159:data<=-32'd473092401;
      160:data<=32'd46078297;
      161:data<=32'd566517123;
      162:data<=32'd1036204963;
      163:data<=32'd1407968501;
      164:data<=32'd1644126095;
      165:data<=32'd1720211545;
      166:data<=32'd1627407330;
      167:data<=32'd1373445063;
      168:data<=32'd981881255;
      169:data<=32'd489816184;
      170:data<=-32'd55723001;
      171:data<=-32'd602381891;
      172:data<=-32'd1097610746;
      173:data<=-32'd1493825108;
      174:data<=-32'd1753087740;
      175:data<=-32'd1850850739;
      176:data<=-32'd1778388378;
      177:data<=-32'd1543679399;
      178:data<=-32'd1170649666;
      179:data<=-32'd696847205;
      180:data<=-32'd169775989;
      181:data<=32'd357752990;
      182:data<=32'd832797646;
      183:data<=32'd1207479648;
      184:data<=32'd1443687609;
      185:data<=32'd1516825814;
      186:data<=32'd1418239018;
      187:data<=32'd1156073616;
      188:data<=32'd754488954;
      189:data<=32'd251294634;
      190:data<=-32'd305755668;
      191:data<=-32'd863651252;
      192:data<=-32'd1369333365;
      193:data<=-32'd1774916137;
      194:data<=-32'd2042409274;
      195:data<=-32'd2147483647;
      196:data<=-32'd2081921335;
      197:data<=-32'd1854539692;
      198:data<=-32'd1490598082;
      199:data<=-32'd1030227337;
      200:data<=-32'd537249431;
      201:data<=32'd55476114;
      202:data<=32'd574438727;
      203:data<=32'd987524279;
      204:data<=32'd1258770772;
      205:data<=32'd1364648650;
      206:data<=32'd1297269858;
      207:data<=32'd1065424378;
      208:data<=32'd693825057;
      209:data<=32'd220735356;
      210:data<=-32'd305755668;
      211:data<=-32'd832432953;
      212:data<=-32'd1306162286;
      213:data<=-32'd1679090247;
      214:data<=-32'd1913325221;
      215:data<=-32'd1984639390;
      216:data<=-32'd1884828446;
      217:data<=-32'd1622498094;
      218:data<=-32'd1222201254;
      219:data<=-32'd722012023;
      220:data<=-32'd169775989;
      221:data<=32'd381593713;
      222:data<=32'd879311847;
      223:data<=32'd1275897483;
      224:data<=32'd1533823312;
      225:data<=32'd1629182189;
      226:data<=32'd1554012351;
      227:data<=32'd1317054992;
      228:data<=32'd942872148;
      229:data<=32'd469414022;
      230:data<=-32'd55723001;
      231:data<=-32'd579978179;
      232:data<=-32'd1050986923;
      233:data<=-32'd1421712643;
      234:data<=-32'd1655046286;
      235:data<=-32'd1727423164;
      236:data<=-32'd1631104030;
      237:data<=-32'd1374899264;
      238:data<=-32'd983268374;
      239:data<=-32'd493886718;
      240:data<=32'd46078297;
      241:data<=32'd584613122;
      242:data<=32'd1069967922;
      243:data<=32'd1455727778;
      244:data<=32'd1705347649;
      245:data<=32'd1795707416;
      246:data<=32'd1719340720;
      247:data<=32'd1485122470;
      248:data<=32'd1117351837;
      249:data<=32'd653325311;
      250:data<=32'd139642436;
      251:data<=-32'd372389462;
      252:data<=-32'd831797781;
      253:data<=-32'd1192938147;
      254:data<=-32'd1419948995;
      255:data<=-32'd1490231849;
      256:data<=-32'd1396619029;
      257:data<=-32'd1148020553;
      258:data<=-32'd768492101;
      259:data<=-32'd294821187;
      260:data<=32'd227126130;
      261:data<=32'd746934815;
      262:data<=32'd1214598782;
      263:data<=32'd1585418943;
      264:data<=32'd1824360864;
      265:data<=32'd1909446559;
      266:data<=32'd1833851526;
      267:data<=32'd1606506677;
      268:data<=32'd1251152556;
      269:data<=32'd803945467;
      270:data<=32'd309857015;
      271:data<=-32'd181774028;
      272:data<=-32'd622096937;
      273:data<=-32'd967532799;
      274:data<=-32'd1184017577;
      275:data<=-32'd1250290611;
      276:data<=-32'd1159910529;
      277:data<=-32'd921807162;
      278:data<=-32'd559322946;
      279:data<=-32'd107845923;
      280:data<=32'd388725618;
      281:data<=32'd882333302;
      282:data<=32'd1325491908;
      283:data<=32'd1675938725;
      284:data<=32'd1900742937;
      285:data<=32'd1979474688;
      286:data<=32'd1906128250;
      287:data<=32'd1689618076;
      288:data<=32'd1352807903;
      289:data<=32'd930177624;
      290:data<=32'd464365906;
      291:data<=32'd1935616;
      292:data<=-32'd411216731;
      293:data<=-32'd734354037;
      294:data<=-32'd935853408;
      295:data<=-32'd996237845;
      296:data<=-32'd909993538;
      297:data<=-32'd686003046;
      298:data<=-32'd346562090;
      299:data<=32'd74912670;
      300:data<=32'd537249431;
      301:data<=32'd995621277;
      302:data<=32'd1405971434;
      303:data<=32'd1729325927;
      304:data<=32'd1935570420;
      305:data<=32'd2006324250;
      306:data<=32'd1936636649;
      307:data<=32'd1735348541;
      308:data<=32'd1424096151;
      309:data<=32'd1035066758;
      310:data<=32'd607738959;
      311:data<=32'd184937884;
      312:data<=-32'd191399715;
      313:data<=-32'd484330602;
      314:data<=-32'd665477365;
      315:data<=-32'd717721292;
      316:data<=-32'd636759482;
      317:data<=-32'd431384542;
      318:data<=-32'd122472877;
      319:data<=32'd259204701;
      320:data<=32'd676121139;
      321:data<=32'd1087759814;
      322:data<=32'd1454630817;
      323:data<=32'd1742137471;
      324:data<=32'd1923913052;
      325:data<=32'd1984304530;
      326:data<=32'd1919768397;
      327:data<=32'd1739054283;
      328:data<=32'd1462173711;
      329:data<=32'd1118271841;
      330:data<=32'd742627451;
      331:data<=32'd373090002;
      332:data<=32'd46314528;
      333:data<=-32'd205829621;
      334:data<=-32'd359322549;
      335:data<=-32'd400233841;
      336:data<=-32'd325928751;
      337:data<=-32'd145136498;
      338:data<=32'd123108399;
      339:data<=32'd451528549;
      340:data<=32'd807448232;
      341:data<=32'd1156123700;
      342:data<=32'd1464218854;
      343:data<=32'd1703076832;
      344:data<=32'd1851464135;
      345:data<=32'd1897522243;
      346:data<=32'd1839745751;
      347:data<=32'd1686907111;
      348:data<=32'd1456955619;
      349:data<=32'd1175021291;
      350:data<=32'd870742391;
      351:data<=32'd575199876;
      352:data<=32'd317776594;
      353:data<=32'd123260801;
      354:data<=32'd9482557;
      355:data<=-32'd14288328;
      356:data<=32'd51963539;
      357:data<=32'd199263280;
      358:data<=32'd410819192;
      359:data<=32'd663963785;
      360:data<=32'd932644335;
      361:data<=32'd1190192353;
      362:data<=32'd1412077905;
      363:data<=32'd1578362297;
      364:data<=32'd1675599984;
      365:data<=32'd1698003401;
      366:data<=32'd1647765751;
      367:data<=32'd1534527889;
      368:data<=32'd1374066483;
      369:data<=32'd1186362086;
      370:data<=32'd993269035;
      371:data<=32'd816047681;
      372:data<=32'd673029448;
      373:data<=32'd577665767;
      374:data<=32'd537165080;
      375:data<=32'd551852609;
      376:data<=32'd615301654;
      377:data<=32'd715188395;
      378:data<=32'd834713313;
      379:data<=32'd954279315;
      380:data<=32'd1052715809;
      381:data<=32'd1104797833;
      382:data<=32'd1064471626;
      383:data<=32'd1070333376;
      384:data<=32'd1076184459;
      385:data<=32'd1082024952;
      386:data<=32'd1087854930;
      387:data<=32'd1093674470;
      388:data<=32'd1099483646;
      389:data<=32'd1105282530;
      390:data<=32'd1111071197;
      391:data<=32'd1116849716;
      392:data<=32'd1122618160;
      393:data<=32'd1128376598;
      394:data<=32'd1134125099;
      395:data<=32'd1139863731;
      396:data<=32'd1145592561;
      397:data<=32'd1151311657;
      398:data<=32'd1157021085;
      399:data<=32'd1162720908;
      400:data<=32'd1168411192;
    endcase
end
assign dout =data;
endmodule
