`timescale 1ns/1ns
package iic_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "iic_transaction.sv"
    `include "iic_sequencer.sv"
    `include "iic_driver.sv"
    `include "iic_monitor.sv"
    `include "iic_agent.sv"
endpackage
